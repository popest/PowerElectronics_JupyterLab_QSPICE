* Coss nonlinear capacitor
.subckt MOS_COSS 1 2
B2 Cp Cn I=V(C_DATA)*DDT(V(Cp,Cn))
R1 2 Cn 1m
R2 1 Cp 1m
B1 C_DATA 0 V=TABLE(abs(V(Cp,Cn)),0,8.75e-09,0.60067,7.69e-09,2.0245,6.63e-09,3.0211,5.74e-09,
+4.8721,4.98e-09,6.723,4.21e-09,9.0418,3.62e-09,11.6352,3.15e-09,16.2625,2.74e-09,
+22.6696,2.46e-09,29.7887,2.29e-09,31.5684,1.95e-09,31.8057,9.84e-10,31.9244,1.7e-09,
+31.9244,1.49e-09,31.9244,1.31e-09,31.9244,1.15e-09,32.0667,3.09e-10,32.2803,5.23e-10,
+32.2803,4.59e-10,32.2803,4.04e-10,32.2803,3.55e-10,32.2803,8.82e-10,32.4939,6.05e-10,
+32.5413,7.44e-10,32.6363,1.97e-10,32.6363,2.71e-10,32.6363,2.38e-10,32.6363,1.62e-10,
+32.6363,1.42e-10,32.7786,7.35e-11,32.9922,1.25e-10,32.9922,1.09e-10,32.9922,9.62e-11,
+32.9922,8.45e-11,33.4905,6.38e-11,34.2635,5.33e-11,36.1958,4.51e-11,38.6366,3.86e-11,
+42.6029,3.34e-11,46.5184,2.95e-11,51.1457,2.61e-11,57.5528,2.29e-11,65.3838,2.05e-11,
+73.2147,1.9e-11,81.0456,1.79e-11,88.8765,1.71e-11,96.7075,1.64e-11,104.5384,1.59e-11,
+112.3693,1.55e-11,120.2002,1.51e-11,128.0311,1.47e-11,135.8621,1.45e-11,143.693,1.42e-11,
+151.5239,1.39e-11,159.3548,1.37e-11,167.1858,1.35e-11,175.0167,1.33e-11,182.8476,1.32e-11,
+190.6785,1.3e-11,198.5095,1.28e-11,206.3404,1.27e-11,214.1713,1.26e-11,222.0022,1.24e-11,
+229.2794,1.23e-11,278.2425,1.17e-11,286.0734,1.16e-11,293.9043,1.16e-11,301.7353,1.15e-11,
+309.5662,1.15e-11,317.3971,1.14e-11,325.228,1.14e-11,333.059,1.13e-11,340.8899,1.13e-11,
+348.7208,1.12e-11,356.5517,1.12e-11,364.3826,1.12e-11,372.2136,1.12e-11,380.0445,1.11e-11,
+387.8754,1.11e-11,395.7063,1.11e-11,403.5373,1.11e-11,411.3682,1.11e-11,419.1991,1.11e-11,
+427.03,1.11e-11,434.861,1.11e-11,442.6919,1.11e-11,450.5228,1.11e-11,458.3537,1.11e-11,
+466.1846,1.11e-11,474.0156,1.11e-11,481.8465,1.11e-11,489.6774,1.11e-11,496.7964,1.11e-11)
.ends MOS_COSS
