* C:\Users\E0481735\OneDrive - Eaton\QSPICE\Input_REC.qsch
D1 N01 out REC
D2 N02 out REC
D3 0 N02 REC
D4 0 N01 REC
V1 N01 N02 SIN 0 {sqrt(2)*VAC_rms} freq
C1 out 0 {Cf}
B1 out 0 R=if(time>1/freq,V(out)*V(out)/{Pin},0)
.model REC D(Vfwd={fwd},Ron={rdiff},Cjo=10p)
.tran 0 {12*1/freq} {1*6/freq} 10�
.options savepowers=1
.param Pin=127.78
.param Cf=116.69�
.param VAC_rms=198
.param fwd=1.2
.param rdiff=0.03
.meas I_AC_RMS rms I(V1)
.meas I_D_RMS rms I(D1)
.meas I_D_AVG avg I(D1)
.meas Pd avg P(V1)
.meas I_Cin_RMS rms I(C1)
.options trtol=1
.meas VOUT_AVG AVG V(out)
.param freq=50
.lib Diode.txt
.end
